// Author: Gong-Chi Wang (王公志)
// NCTU IC Lab Exercise #1
//================================================================
//   File Name   : sort.v
//   Module Name : Sort
//   Description : Sort the input signals (ID/Gm) in ascending order, *with combination logic only, i.e., no clk*
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

module Sort(
    // Input signals
    in0, in1, in2, in3, in4, in5,
    mode,
    // Output signals
    out0, out1, out2, out3, out4, out5
);
input [6:0] in0, in1, in2, in3, in4, in5;
input mode; // 0: Ascending, 1: Descending
output [6:0] out0, out1, out2, out3, out4, out5;





endmodule
